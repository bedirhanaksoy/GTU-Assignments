module move(output [31:0] moved_rt, input [31:0] rs);

  and and1(moved_rt[0], rs[0], 1'b1);
  and and2(moved_rt[1], rs[1], 1'b1);
  and and3(moved_rt[2], rs[2], 1'b1);
  and and4(moved_rt[3], rs[3], 1'b1);
  and and5(moved_rt[4], rs[4], 1'b1);
  and and6(moved_rt[5], rs[5], 1'b1);
  and and7(moved_rt[6], rs[6], 1'b1);
  and and8(moved_rt[7], rs[7], 1'b1);
  and and9(moved_rt[8], rs[8], 1'b1);
  and and10(moved_rt[9], rs[9], 1'b1);
  and and11(moved_rt[10], rs[10], 1'b1);
  and and12(moved_rt[11], rs[11], 1'b1);
  and and13(moved_rt[12], rs[12], 1'b1);
  and and14(moved_rt[13], rs[13], 1'b1);
  and and15(moved_rt[14], rs[14], 1'b1);
  and and16(moved_rt[15], rs[15], 1'b1);
  and and17(moved_rt[16], rs[16], 1'b1);
  and and18(moved_rt[17], rs[17], 1'b1);
  and and19(moved_rt[18], rs[18], 1'b1);
  and and20(moved_rt[19], rs[19], 1'b1);
  and and21(moved_rt[20], rs[20], 1'b1);
  and and22(moved_rt[21], rs[21], 1'b1);
  and and23(moved_rt[22], rs[22], 1'b1);
  and and24(moved_rt[23], rs[23], 1'b1);
  and and25(moved_rt[24], rs[24], 1'b1);
  and and26(moved_rt[25], rs[25], 1'b1);
  and and27(moved_rt[26], rs[26], 1'b1);
  and and28(moved_rt[27], rs[27], 1'b1);
  and and29(moved_rt[28], rs[28], 1'b1);
  and and30(moved_rt[29], rs[29], 1'b1);
  and and31(moved_rt[30], rs[30], 1'b1);
  and and32(moved_rt[31], rs[31], 1'b1);

endmodule
