module PC_four_adder(input [31:0] PC, output [31:0] incremented_PC);

thirty_two_bit_adder(

endmodule
