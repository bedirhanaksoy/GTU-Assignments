module PC_mux(input [31:0] PC_4_add_result, 
				  input [31:0] PC_shift_left_add_result, 
				  input zero_and_branch, 
				  output [31:0] PC);

  wire [31:0] temp_res1;
  wire [31:0] temp_res2;
  wire zero_and_branch_;

  not not1(zero_and_branch_, zero_and_branch);

  and and1(temp_res1[31], PC_4_add_result[31], zero_and_branch_);
  and and2(temp_res1[30], PC_4_add_result[30], zero_and_branch_);
  and and3(temp_res1[29], PC_4_add_result[29], zero_and_branch_);
  and and4(temp_res1[28], PC_4_add_result[28], zero_and_branch_);
  and and5(temp_res1[27], PC_4_add_result[27], zero_and_branch_);
  and and6(temp_res1[26], PC_4_add_result[26], zero_and_branch_);
  and and7(temp_res1[25], PC_4_add_result[25], zero_and_branch_);
  and and8(temp_res1[24], PC_4_add_result[24], zero_and_branch_);
  and and9(temp_res1[23], PC_4_add_result[23], zero_and_branch_);
  and and10(temp_res1[22], PC_4_add_result[22], zero_and_branch_);
  and and11(temp_res1[21], PC_4_add_result[21], zero_and_branch_);
  and and12(temp_res1[20], PC_4_add_result[20], zero_and_branch_);
  and and13(temp_res1[19], PC_4_add_result[19], zero_and_branch_);
  and and14(temp_res1[18], PC_4_add_result[18], zero_and_branch_);
  and and15(temp_res1[17], PC_4_add_result[17], zero_and_branch_);
  and and16(temp_res1[16], PC_4_add_result[16], zero_and_branch_);
  and and17(temp_res1[15], PC_4_add_result[15], zero_and_branch_);
  and and18(temp_res1[14], PC_4_add_result[14], zero_and_branch_);
  and and19(temp_res1[13], PC_4_add_result[13], zero_and_branch_);
  and and20(temp_res1[12], PC_4_add_result[12], zero_and_branch_);
  and and21(temp_res1[11], PC_4_add_result[11], zero_and_branch_);
  and and22(temp_res1[10], PC_4_add_result[10], zero_and_branch_);
  and and23(temp_res1[9], PC_4_add_result[9], zero_and_branch_);
  and and24(temp_res1[8], PC_4_add_result[8], zero_and_branch_);
  and and25(temp_res1[7], PC_4_add_result[7], zero_and_branch_);
  and and26(temp_res1[6], PC_4_add_result[6], zero_and_branch_);
  and and27(temp_res1[5], PC_4_add_result[5], zero_and_branch_);
  and and28(temp_res1[4], PC_4_add_result[4], zero_and_branch_);
  and and29(temp_res1[3], PC_4_add_result[3], zero_and_branch_);
  and and30(temp_res1[2], PC_4_add_result[2], zero_and_branch_);
  and and31(temp_res1[1], PC_4_add_result[1], zero_and_branch_);
  and and32(temp_res1[0], PC_4_add_result[0], zero_and_branch_);

  and and33(temp_res2[31], PC_shift_left_add_result[31], zero_and_branch);
  and and34(temp_res2[30], PC_shift_left_add_result[30], zero_and_branch);
  and and35(temp_res2[29], PC_shift_left_add_result[29], zero_and_branch);
  and and36(temp_res2[28], PC_shift_left_add_result[28], zero_and_branch);
  and and37(temp_res2[27], PC_shift_left_add_result[27], zero_and_branch);
  and and38(temp_res2[26], PC_shift_left_add_result[26], zero_and_branch);
  and and39(temp_res2[25], PC_shift_left_add_result[25], zero_and_branch);
  and and40(temp_res2[24], PC_shift_left_add_result[24], zero_and_branch);
  and and41(temp_res2[23], PC_shift_left_add_result[23], zero_and_branch);
  and and42(temp_res2[22], PC_shift_left_add_result[22], zero_and_branch);
  and and43(temp_res2[21], PC_shift_left_add_result[21], zero_and_branch);
  and and44(temp_res2[20], PC_shift_left_add_result[20], zero_and_branch);
  and and45(temp_res2[19], PC_shift_left_add_result[19], zero_and_branch);
  and and46(temp_res2[18], PC_shift_left_add_result[18], zero_and_branch);
  and and47(temp_res2[17], PC_shift_left_add_result[17], zero_and_branch);
  and and48(temp_res2[16], PC_shift_left_add_result[16], zero_and_branch);
  and and49(temp_res2[15], PC_shift_left_add_result[15], zero_and_branch);
  and and50(temp_res2[14], PC_shift_left_add_result[14], zero_and_branch);
  and and51(temp_res2[13], PC_shift_left_add_result[13], zero_and_branch);
  and and52(temp_res2[12], PC_shift_left_add_result[12], zero_and_branch);
  and and53(temp_res2[11], PC_shift_left_add_result[11], zero_and_branch);
  and and54(temp_res2[10], PC_shift_left_add_result[10], zero_and_branch);
  and and55(temp_res2[9], PC_shift_left_add_result[9], zero_and_branch);
  and and56(temp_res2[8], PC_shift_left_add_result[8], zero_and_branch);
  and and57(temp_res2[7], PC_shift_left_add_result[7], zero_and_branch);
  and and58(temp_res2[6], PC_shift_left_add_result[6], zero_and_branch);
  and and59(temp_res2[5], PC_shift_left_add_result[5], zero_and_branch);
  and and60(temp_res2[4], PC_shift_left_add_result[4], zero_and_branch);
  and and61(temp_res2[3], PC_shift_left_add_result[3], zero_and_branch);
  and and62(temp_res2[2], PC_shift_left_add_result[2], zero_and_branch);
  and and63(temp_res2[1], PC_shift_left_add_result[1], zero_and_branch);
  and and64(temp_res2[0], PC_shift_left_add_result[0], zero_and_branch);

  or or1(PC[31], temp_res1[31], temp_res2[31]);
  or or2(PC[30], temp_res1[30], temp_res2[30]);
  or or3(PC[29], temp_res1[29], temp_res2[29]);
  or or4(PC[28], temp_res1[28], temp_res2[28]);
  or or5(PC[27], temp_res1[27], temp_res2[27]);
  or or6(PC[26], temp_res1[26], temp_res2[26]);
  or or7(PC[25], temp_res1[25], temp_res2[25]);
  or or8(PC[24], temp_res1[24], temp_res2[24]);
  or or9(PC[23], temp_res1[23], temp_res2[23]);
  or or10(PC[22], temp_res1[22], temp_res2[22]);
  or or11(PC[21], temp_res1[21], temp_res2[21]);
  or or12(PC[20], temp_res1[20], temp_res2[20]);
  or or13(PC[19], temp_res1[19], temp_res2[19]);
  or or14(PC[18], temp_res1[18], temp_res2[18]);
  or or15(PC[17], temp_res1[17], temp_res2[17]);
  or or16(PC[16], temp_res1[16], temp_res2[16]);
  or or17(PC[15], temp_res1[15], temp_res2[15]);
  or or18(PC[14], temp_res1[14], temp_res2[14]);
  or or19(PC[13], temp_res1[13], temp_res2[13]);
  or or20(PC[12], temp_res1[12], temp_res2[12]);
  or or21(PC[11], temp_res1[11], temp_res2[11]);
  or or22(PC[10], temp_res1[10], temp_res2[10]);
  or or23(PC[9], temp_res1[9], temp_res2[9]);
  or or24(PC[8], temp_res1[8], temp_res2[8]);
  or or25(PC[7], temp_res1[7], temp_res2[7]);
  or or26(PC[6], temp_res1[6], temp_res2[6]);
  or or27(PC[5], temp_res1[5], temp_res2[5]);
  or or28(PC[4], temp_res1[4], temp_res2[4]);
  or or29(PC[3], temp_res1[3], temp_res2[3]);
  or or30(PC[2], temp_res1[2], temp_res2[2]);
  or or31(PC[1], temp_res1[1], temp_res2[1]);
  or or32(PC[0], temp_res1[0], temp_res2[0]);

endmodule
