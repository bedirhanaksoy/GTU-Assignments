module mipstestbench(input clk);

mips test1(clk);

endmodule
